
module mem_MM #(                   // 
    parameter  ADDR_LEN  = 11   // 
) (
    input  clk, rst,
    input  [ADDR_LEN-1:0] addr, // memory address
    output reg [31:0] rd_data,  // data read out
    input  wr_req,
    input  [31:0] wr_data       // data write in
);
localparam MEM_SIZE = 1<<ADDR_LEN;
reg [31:0] ram_cell [MEM_SIZE];

always @ (posedge clk or posedge rst)
    if(rst)
        rd_data <= 0;
    else
        rd_data <= ram_cell[addr];

always @ (posedge clk)
    if(wr_req) 
        ram_cell[addr] <= wr_data;

initial begin
    // dst matrix C
    ram_cell[       0] = 32'h0;  // 32'h318e4a02;
    ram_cell[       1] = 32'h0;  // 32'hb9c70164;
    ram_cell[       2] = 32'h0;  // 32'h1b1d6c1d;
    ram_cell[       3] = 32'h0;  // 32'h6cf187a3;
    ram_cell[       4] = 32'h0;  // 32'h3312eced;
    ram_cell[       5] = 32'h0;  // 32'he1f6b8c8;
    ram_cell[       6] = 32'h0;  // 32'h042c1a66;
    ram_cell[       7] = 32'h0;  // 32'h52238a15;
    ram_cell[       8] = 32'h0;  // 32'hcee8d2ab;
    ram_cell[       9] = 32'h0;  // 32'h60c9fe6b;
    ram_cell[      10] = 32'h0;  // 32'h919d7d8f;
    ram_cell[      11] = 32'h0;  // 32'h6b62a2f3;
    ram_cell[      12] = 32'h0;  // 32'hc848704c;
    ram_cell[      13] = 32'h0;  // 32'h3a88c347;
    ram_cell[      14] = 32'h0;  // 32'h4745ef41;
    ram_cell[      15] = 32'h0;  // 32'h9cde7860;
    ram_cell[      16] = 32'h0;  // 32'hbc56972b;
    ram_cell[      17] = 32'h0;  // 32'hd33aad10;
    ram_cell[      18] = 32'h0;  // 32'h3a71c723;
    ram_cell[      19] = 32'h0;  // 32'h6a72054c;
    ram_cell[      20] = 32'h0;  // 32'hc387c2a0;
    ram_cell[      21] = 32'h0;  // 32'h492375e0;
    ram_cell[      22] = 32'h0;  // 32'hd98caf78;
    ram_cell[      23] = 32'h0;  // 32'h6f3830ba;
    ram_cell[      24] = 32'h0;  // 32'hed50c911;
    ram_cell[      25] = 32'h0;  // 32'h84c47c38;
    ram_cell[      26] = 32'h0;  // 32'h6f517d6b;
    ram_cell[      27] = 32'h0;  // 32'ha2b93106;
    ram_cell[      28] = 32'h0;  // 32'h47fadbaf;
    ram_cell[      29] = 32'h0;  // 32'h0ed0a615;
    ram_cell[      30] = 32'h0;  // 32'h1dc1893f;
    ram_cell[      31] = 32'h0;  // 32'h9db04777;
    ram_cell[      32] = 32'h0;  // 32'h39683d09;
    ram_cell[      33] = 32'h0;  // 32'h779d038d;
    ram_cell[      34] = 32'h0;  // 32'h726a0b3e;
    ram_cell[      35] = 32'h0;  // 32'hb3e9bb3f;
    ram_cell[      36] = 32'h0;  // 32'h3268d31e;
    ram_cell[      37] = 32'h0;  // 32'h3f1aeb68;
    ram_cell[      38] = 32'h0;  // 32'hfc2804de;
    ram_cell[      39] = 32'h0;  // 32'h8382c4e1;
    ram_cell[      40] = 32'h0;  // 32'h8b714ba1;
    ram_cell[      41] = 32'h0;  // 32'hfd7b264c;
    ram_cell[      42] = 32'h0;  // 32'hc6931a40;
    ram_cell[      43] = 32'h0;  // 32'h60a77571;
    ram_cell[      44] = 32'h0;  // 32'hcb3a7ce8;
    ram_cell[      45] = 32'h0;  // 32'h0de0267e;
    ram_cell[      46] = 32'h0;  // 32'h02b85e71;
    ram_cell[      47] = 32'h0;  // 32'ha34c46c3;
    ram_cell[      48] = 32'h0;  // 32'h9bca6677;
    ram_cell[      49] = 32'h0;  // 32'h925c5fb5;
    ram_cell[      50] = 32'h0;  // 32'hdfd35146;
    ram_cell[      51] = 32'h0;  // 32'h28747560;
    ram_cell[      52] = 32'h0;  // 32'h90bd6da5;
    ram_cell[      53] = 32'h0;  // 32'h7e0091a8;
    ram_cell[      54] = 32'h0;  // 32'h148d90ce;
    ram_cell[      55] = 32'h0;  // 32'h1a8f0954;
    ram_cell[      56] = 32'h0;  // 32'hecffc05d;
    ram_cell[      57] = 32'h0;  // 32'hec46e588;
    ram_cell[      58] = 32'h0;  // 32'h1d2d4108;
    ram_cell[      59] = 32'h0;  // 32'hf7412209;
    ram_cell[      60] = 32'h0;  // 32'h4dbe546b;
    ram_cell[      61] = 32'h0;  // 32'h4831727a;
    ram_cell[      62] = 32'h0;  // 32'h267389bb;
    ram_cell[      63] = 32'h0;  // 32'h92118284;
    ram_cell[      64] = 32'h0;  // 32'h56e4217f;
    ram_cell[      65] = 32'h0;  // 32'h780d0f66;
    ram_cell[      66] = 32'h0;  // 32'h6ddb780a;
    ram_cell[      67] = 32'h0;  // 32'hd83fbe1b;
    ram_cell[      68] = 32'h0;  // 32'h036f5e0b;
    ram_cell[      69] = 32'h0;  // 32'h06a5cb24;
    ram_cell[      70] = 32'h0;  // 32'h49182db6;
    ram_cell[      71] = 32'h0;  // 32'h40f7d573;
    ram_cell[      72] = 32'h0;  // 32'h6f7ea02d;
    ram_cell[      73] = 32'h0;  // 32'h13846e55;
    ram_cell[      74] = 32'h0;  // 32'h1c3ec10c;
    ram_cell[      75] = 32'h0;  // 32'h53cdba88;
    ram_cell[      76] = 32'h0;  // 32'he88952c1;
    ram_cell[      77] = 32'h0;  // 32'h95f0e7dc;
    ram_cell[      78] = 32'h0;  // 32'h019ff2c4;
    ram_cell[      79] = 32'h0;  // 32'h54458530;
    ram_cell[      80] = 32'h0;  // 32'h5f355cdd;
    ram_cell[      81] = 32'h0;  // 32'h493c75ff;
    ram_cell[      82] = 32'h0;  // 32'h0e937c93;
    ram_cell[      83] = 32'h0;  // 32'h54200fd6;
    ram_cell[      84] = 32'h0;  // 32'hd0adeb41;
    ram_cell[      85] = 32'h0;  // 32'h434c9199;
    ram_cell[      86] = 32'h0;  // 32'hd289e435;
    ram_cell[      87] = 32'h0;  // 32'hd2ed15d3;
    ram_cell[      88] = 32'h0;  // 32'ha05faf56;
    ram_cell[      89] = 32'h0;  // 32'ha20b92c5;
    ram_cell[      90] = 32'h0;  // 32'hc9e92a6d;
    ram_cell[      91] = 32'h0;  // 32'h9cc58b9a;
    ram_cell[      92] = 32'h0;  // 32'h27f83eb0;
    ram_cell[      93] = 32'h0;  // 32'h03b931ef;
    ram_cell[      94] = 32'h0;  // 32'h01a2ad15;
    ram_cell[      95] = 32'h0;  // 32'h12b1bf41;
    ram_cell[      96] = 32'h0;  // 32'h37e97031;
    ram_cell[      97] = 32'h0;  // 32'h3c64c58d;
    ram_cell[      98] = 32'h0;  // 32'h1a3aef68;
    ram_cell[      99] = 32'h0;  // 32'h5520931c;
    ram_cell[     100] = 32'h0;  // 32'h3fce8b2b;
    ram_cell[     101] = 32'h0;  // 32'hae45abf6;
    ram_cell[     102] = 32'h0;  // 32'h50de8ef7;
    ram_cell[     103] = 32'h0;  // 32'h2cea9c6a;
    ram_cell[     104] = 32'h0;  // 32'h23719ba3;
    ram_cell[     105] = 32'h0;  // 32'hc22bde11;
    ram_cell[     106] = 32'h0;  // 32'h97ffa26d;
    ram_cell[     107] = 32'h0;  // 32'h3cc0f182;
    ram_cell[     108] = 32'h0;  // 32'h49e7c5f4;
    ram_cell[     109] = 32'h0;  // 32'h83698b6c;
    ram_cell[     110] = 32'h0;  // 32'hf5e4666a;
    ram_cell[     111] = 32'h0;  // 32'hfd3b79b8;
    ram_cell[     112] = 32'h0;  // 32'h3ea2261f;
    ram_cell[     113] = 32'h0;  // 32'h30fcb009;
    ram_cell[     114] = 32'h0;  // 32'h771960ff;
    ram_cell[     115] = 32'h0;  // 32'h3db8ad42;
    ram_cell[     116] = 32'h0;  // 32'h796cbedf;
    ram_cell[     117] = 32'h0;  // 32'h9f17662a;
    ram_cell[     118] = 32'h0;  // 32'hc11cea3b;
    ram_cell[     119] = 32'h0;  // 32'h3560b0bd;
    ram_cell[     120] = 32'h0;  // 32'h2304654f;
    ram_cell[     121] = 32'h0;  // 32'hf79428bd;
    ram_cell[     122] = 32'h0;  // 32'h83c31eac;
    ram_cell[     123] = 32'h0;  // 32'hd939a802;
    ram_cell[     124] = 32'h0;  // 32'hc6b3099d;
    ram_cell[     125] = 32'h0;  // 32'hac204fc6;
    ram_cell[     126] = 32'h0;  // 32'h5b155311;
    ram_cell[     127] = 32'h0;  // 32'h0c6334f6;
    ram_cell[     128] = 32'h0;  // 32'h2e17be7b;
    ram_cell[     129] = 32'h0;  // 32'h0cf6c068;
    ram_cell[     130] = 32'h0;  // 32'h7fc2562f;
    ram_cell[     131] = 32'h0;  // 32'h44d19d3f;
    ram_cell[     132] = 32'h0;  // 32'h029b7f9b;
    ram_cell[     133] = 32'h0;  // 32'hb8f80eb5;
    ram_cell[     134] = 32'h0;  // 32'h7fb72af3;
    ram_cell[     135] = 32'h0;  // 32'h2a1408bb;
    ram_cell[     136] = 32'h0;  // 32'h8170bd99;
    ram_cell[     137] = 32'h0;  // 32'ha98a8d01;
    ram_cell[     138] = 32'h0;  // 32'h7da68b9f;
    ram_cell[     139] = 32'h0;  // 32'h2ae9eb61;
    ram_cell[     140] = 32'h0;  // 32'h05efa847;
    ram_cell[     141] = 32'h0;  // 32'hfc48d794;
    ram_cell[     142] = 32'h0;  // 32'hcb2643d4;
    ram_cell[     143] = 32'h0;  // 32'hcde2e0e3;
    ram_cell[     144] = 32'h0;  // 32'h7fa0d83f;
    ram_cell[     145] = 32'h0;  // 32'h8ef74552;
    ram_cell[     146] = 32'h0;  // 32'he1702ed3;
    ram_cell[     147] = 32'h0;  // 32'h5c9d556f;
    ram_cell[     148] = 32'h0;  // 32'h192e2444;
    ram_cell[     149] = 32'h0;  // 32'ha8d00ace;
    ram_cell[     150] = 32'h0;  // 32'h4d37b9eb;
    ram_cell[     151] = 32'h0;  // 32'haf762125;
    ram_cell[     152] = 32'h0;  // 32'ha7214de4;
    ram_cell[     153] = 32'h0;  // 32'h3d3e668e;
    ram_cell[     154] = 32'h0;  // 32'h8edb689c;
    ram_cell[     155] = 32'h0;  // 32'h1e2badcb;
    ram_cell[     156] = 32'h0;  // 32'h6782db24;
    ram_cell[     157] = 32'h0;  // 32'h28343e41;
    ram_cell[     158] = 32'h0;  // 32'h7a60e530;
    ram_cell[     159] = 32'h0;  // 32'ha5db9e46;
    ram_cell[     160] = 32'h0;  // 32'h579d5dbe;
    ram_cell[     161] = 32'h0;  // 32'hb71e792b;
    ram_cell[     162] = 32'h0;  // 32'he12e553e;
    ram_cell[     163] = 32'h0;  // 32'h44d504c5;
    ram_cell[     164] = 32'h0;  // 32'hd6b5fd78;
    ram_cell[     165] = 32'h0;  // 32'h350e1754;
    ram_cell[     166] = 32'h0;  // 32'h4eba73fa;
    ram_cell[     167] = 32'h0;  // 32'hd2707d0e;
    ram_cell[     168] = 32'h0;  // 32'h819f9469;
    ram_cell[     169] = 32'h0;  // 32'h184ec423;
    ram_cell[     170] = 32'h0;  // 32'h5da554d3;
    ram_cell[     171] = 32'h0;  // 32'h5a5fdf65;
    ram_cell[     172] = 32'h0;  // 32'hbe03871b;
    ram_cell[     173] = 32'h0;  // 32'h91443f4b;
    ram_cell[     174] = 32'h0;  // 32'hcf69f28a;
    ram_cell[     175] = 32'h0;  // 32'h2f59810f;
    ram_cell[     176] = 32'h0;  // 32'h8a65d82f;
    ram_cell[     177] = 32'h0;  // 32'h20f7989f;
    ram_cell[     178] = 32'h0;  // 32'h71b10f7f;
    ram_cell[     179] = 32'h0;  // 32'h54dd5db3;
    ram_cell[     180] = 32'h0;  // 32'haf21566a;
    ram_cell[     181] = 32'h0;  // 32'h7a5ec1af;
    ram_cell[     182] = 32'h0;  // 32'he54a8598;
    ram_cell[     183] = 32'h0;  // 32'h11f11e17;
    ram_cell[     184] = 32'h0;  // 32'hc8e167a8;
    ram_cell[     185] = 32'h0;  // 32'h065e5f50;
    ram_cell[     186] = 32'h0;  // 32'h1993eca3;
    ram_cell[     187] = 32'h0;  // 32'h73d11555;
    ram_cell[     188] = 32'h0;  // 32'ha5a2c0d9;
    ram_cell[     189] = 32'h0;  // 32'h2f65fa04;
    ram_cell[     190] = 32'h0;  // 32'hce975b4b;
    ram_cell[     191] = 32'h0;  // 32'hceadd778;
    ram_cell[     192] = 32'h0;  // 32'h9560ccb8;
    ram_cell[     193] = 32'h0;  // 32'hb875a086;
    ram_cell[     194] = 32'h0;  // 32'h8b65b4b6;
    ram_cell[     195] = 32'h0;  // 32'h5fb8dfde;
    ram_cell[     196] = 32'h0;  // 32'hd8d41c34;
    ram_cell[     197] = 32'h0;  // 32'hb480ed1e;
    ram_cell[     198] = 32'h0;  // 32'hc9217e23;
    ram_cell[     199] = 32'h0;  // 32'h5e6dad56;
    ram_cell[     200] = 32'h0;  // 32'h325294b4;
    ram_cell[     201] = 32'h0;  // 32'h768bdbd4;
    ram_cell[     202] = 32'h0;  // 32'haca3eddd;
    ram_cell[     203] = 32'h0;  // 32'h7c0cb53e;
    ram_cell[     204] = 32'h0;  // 32'hf393c26c;
    ram_cell[     205] = 32'h0;  // 32'h5482e817;
    ram_cell[     206] = 32'h0;  // 32'hd03c2c4c;
    ram_cell[     207] = 32'h0;  // 32'hc840c531;
    ram_cell[     208] = 32'h0;  // 32'hb21be36b;
    ram_cell[     209] = 32'h0;  // 32'h2da67ec2;
    ram_cell[     210] = 32'h0;  // 32'h96936d30;
    ram_cell[     211] = 32'h0;  // 32'h60d94ebd;
    ram_cell[     212] = 32'h0;  // 32'h779823ba;
    ram_cell[     213] = 32'h0;  // 32'hb14e8ec4;
    ram_cell[     214] = 32'h0;  // 32'h8af7f327;
    ram_cell[     215] = 32'h0;  // 32'h3b206744;
    ram_cell[     216] = 32'h0;  // 32'h88abdf80;
    ram_cell[     217] = 32'h0;  // 32'ha0cbb2af;
    ram_cell[     218] = 32'h0;  // 32'h9c730703;
    ram_cell[     219] = 32'h0;  // 32'h22aaa7a0;
    ram_cell[     220] = 32'h0;  // 32'hb02d4432;
    ram_cell[     221] = 32'h0;  // 32'h5d356b15;
    ram_cell[     222] = 32'h0;  // 32'h0d5926d8;
    ram_cell[     223] = 32'h0;  // 32'h8fe3fb43;
    ram_cell[     224] = 32'h0;  // 32'h3269e7e6;
    ram_cell[     225] = 32'h0;  // 32'h168f88ec;
    ram_cell[     226] = 32'h0;  // 32'h8ea5e171;
    ram_cell[     227] = 32'h0;  // 32'hb54e8177;
    ram_cell[     228] = 32'h0;  // 32'h77f3dd8e;
    ram_cell[     229] = 32'h0;  // 32'h3b3f7285;
    ram_cell[     230] = 32'h0;  // 32'h04904125;
    ram_cell[     231] = 32'h0;  // 32'h900d701d;
    ram_cell[     232] = 32'h0;  // 32'hdc65f8a2;
    ram_cell[     233] = 32'h0;  // 32'h4f3ab136;
    ram_cell[     234] = 32'h0;  // 32'he533539f;
    ram_cell[     235] = 32'h0;  // 32'h13665185;
    ram_cell[     236] = 32'h0;  // 32'hf1750065;
    ram_cell[     237] = 32'h0;  // 32'h80270321;
    ram_cell[     238] = 32'h0;  // 32'h4223a902;
    ram_cell[     239] = 32'h0;  // 32'h306703a6;
    ram_cell[     240] = 32'h0;  // 32'h8f6edee9;
    ram_cell[     241] = 32'h0;  // 32'h011b58f3;
    ram_cell[     242] = 32'h0;  // 32'h9be14098;
    ram_cell[     243] = 32'h0;  // 32'ha486dc0b;
    ram_cell[     244] = 32'h0;  // 32'h4248319a;
    ram_cell[     245] = 32'h0;  // 32'h3db2bca2;
    ram_cell[     246] = 32'h0;  // 32'hb172e506;
    ram_cell[     247] = 32'h0;  // 32'hc810334f;
    ram_cell[     248] = 32'h0;  // 32'h6f1d3478;
    ram_cell[     249] = 32'h0;  // 32'h5fb6488b;
    ram_cell[     250] = 32'h0;  // 32'hd32d65c4;
    ram_cell[     251] = 32'h0;  // 32'h7e1553bc;
    ram_cell[     252] = 32'h0;  // 32'h80d6b2bf;
    ram_cell[     253] = 32'h0;  // 32'hd4c6a848;
    ram_cell[     254] = 32'h0;  // 32'h4932dc57;
    ram_cell[     255] = 32'h0;  // 32'h4f09a056;
    // src matrix A
    ram_cell[     256] = 32'h00dd6be0;
    ram_cell[     257] = 32'h42cbce48;
    ram_cell[     258] = 32'hc78fe644;
    ram_cell[     259] = 32'hdcc93307;
    ram_cell[     260] = 32'heb158c89;
    ram_cell[     261] = 32'hc0dabf5c;
    ram_cell[     262] = 32'h25a79ede;
    ram_cell[     263] = 32'hb16f2b0f;
    ram_cell[     264] = 32'h4d4dfa1f;
    ram_cell[     265] = 32'h8881f864;
    ram_cell[     266] = 32'h76a78561;
    ram_cell[     267] = 32'hfcff9ecb;
    ram_cell[     268] = 32'h7f4dbfd3;
    ram_cell[     269] = 32'haedccc4a;
    ram_cell[     270] = 32'he73b2f4a;
    ram_cell[     271] = 32'h4d37f20e;
    ram_cell[     272] = 32'hec4f7eea;
    ram_cell[     273] = 32'h21c03f7b;
    ram_cell[     274] = 32'h336b894f;
    ram_cell[     275] = 32'h14201bc5;
    ram_cell[     276] = 32'h4c65992a;
    ram_cell[     277] = 32'h7a5a6c97;
    ram_cell[     278] = 32'h8d0ead8e;
    ram_cell[     279] = 32'h6a4ce672;
    ram_cell[     280] = 32'h4cce6b40;
    ram_cell[     281] = 32'hd4d8cf15;
    ram_cell[     282] = 32'ha3954320;
    ram_cell[     283] = 32'h7a659c9e;
    ram_cell[     284] = 32'h7a9a2d0c;
    ram_cell[     285] = 32'hce199294;
    ram_cell[     286] = 32'h023e87b5;
    ram_cell[     287] = 32'h4e5512dc;
    ram_cell[     288] = 32'hecd0278f;
    ram_cell[     289] = 32'he150b98c;
    ram_cell[     290] = 32'ha0a8b2bc;
    ram_cell[     291] = 32'he0875fc7;
    ram_cell[     292] = 32'hcf193c52;
    ram_cell[     293] = 32'hf04f5c03;
    ram_cell[     294] = 32'h546433cc;
    ram_cell[     295] = 32'hd4bfbca2;
    ram_cell[     296] = 32'hc5695161;
    ram_cell[     297] = 32'h79028f8a;
    ram_cell[     298] = 32'h42a33cc3;
    ram_cell[     299] = 32'hd5d6d525;
    ram_cell[     300] = 32'h22108326;
    ram_cell[     301] = 32'h9bcc886b;
    ram_cell[     302] = 32'h57ba950d;
    ram_cell[     303] = 32'hda07359f;
    ram_cell[     304] = 32'hf80e6699;
    ram_cell[     305] = 32'h149aa21b;
    ram_cell[     306] = 32'h993d6874;
    ram_cell[     307] = 32'h19f9ebb3;
    ram_cell[     308] = 32'h1fbb3540;
    ram_cell[     309] = 32'h193ab402;
    ram_cell[     310] = 32'h63afd5b6;
    ram_cell[     311] = 32'h0e4368aa;
    ram_cell[     312] = 32'h1245beed;
    ram_cell[     313] = 32'h1991c42f;
    ram_cell[     314] = 32'hb0f3d81d;
    ram_cell[     315] = 32'h4fa072fe;
    ram_cell[     316] = 32'h83fb0f48;
    ram_cell[     317] = 32'h89979a52;
    ram_cell[     318] = 32'h69451c2d;
    ram_cell[     319] = 32'hb2051155;
    ram_cell[     320] = 32'h498e06dd;
    ram_cell[     321] = 32'h0b7e6eff;
    ram_cell[     322] = 32'h546b5db5;
    ram_cell[     323] = 32'h24d21433;
    ram_cell[     324] = 32'hc82129a8;
    ram_cell[     325] = 32'h74975d29;
    ram_cell[     326] = 32'h1d85d469;
    ram_cell[     327] = 32'h146feb75;
    ram_cell[     328] = 32'h12c5bfe1;
    ram_cell[     329] = 32'hcb48fe92;
    ram_cell[     330] = 32'h0f9a8414;
    ram_cell[     331] = 32'he748fca0;
    ram_cell[     332] = 32'h05d77fab;
    ram_cell[     333] = 32'h2f03859f;
    ram_cell[     334] = 32'h2f5e9f3d;
    ram_cell[     335] = 32'h2f9e5b17;
    ram_cell[     336] = 32'h98a4a49b;
    ram_cell[     337] = 32'h4fbd8256;
    ram_cell[     338] = 32'h81ed53e9;
    ram_cell[     339] = 32'he241d270;
    ram_cell[     340] = 32'hd4a89cc0;
    ram_cell[     341] = 32'h9a7d147c;
    ram_cell[     342] = 32'h4dbbee25;
    ram_cell[     343] = 32'h008146d2;
    ram_cell[     344] = 32'h1f73bfa8;
    ram_cell[     345] = 32'h01221a0b;
    ram_cell[     346] = 32'h31402f50;
    ram_cell[     347] = 32'h5df765b1;
    ram_cell[     348] = 32'h67851fc1;
    ram_cell[     349] = 32'hb32ee917;
    ram_cell[     350] = 32'ha0cf2f6e;
    ram_cell[     351] = 32'h7c88c462;
    ram_cell[     352] = 32'h0c260c8d;
    ram_cell[     353] = 32'hddd6814f;
    ram_cell[     354] = 32'h6bc2c458;
    ram_cell[     355] = 32'h87e31435;
    ram_cell[     356] = 32'h1b3241ff;
    ram_cell[     357] = 32'he5b50fa1;
    ram_cell[     358] = 32'h1c146f9f;
    ram_cell[     359] = 32'h3f656aa2;
    ram_cell[     360] = 32'h6baaafc8;
    ram_cell[     361] = 32'h1cee20d6;
    ram_cell[     362] = 32'h5c75ccb0;
    ram_cell[     363] = 32'hb5e72f2e;
    ram_cell[     364] = 32'h59077262;
    ram_cell[     365] = 32'hdc262724;
    ram_cell[     366] = 32'h8c6b133e;
    ram_cell[     367] = 32'h1e38dfa1;
    ram_cell[     368] = 32'h0d1fcb8c;
    ram_cell[     369] = 32'h395ed167;
    ram_cell[     370] = 32'h80c39ae1;
    ram_cell[     371] = 32'hc4ddee4a;
    ram_cell[     372] = 32'h955c9b73;
    ram_cell[     373] = 32'hf63e90a2;
    ram_cell[     374] = 32'h1381a51a;
    ram_cell[     375] = 32'h744785c8;
    ram_cell[     376] = 32'he893aeaa;
    ram_cell[     377] = 32'h2c3463a9;
    ram_cell[     378] = 32'h654cbd63;
    ram_cell[     379] = 32'hf2227a61;
    ram_cell[     380] = 32'h047782ff;
    ram_cell[     381] = 32'h31e79934;
    ram_cell[     382] = 32'hdc3cc4b8;
    ram_cell[     383] = 32'hd1081bb9;
    ram_cell[     384] = 32'h9cd1fbf7;
    ram_cell[     385] = 32'h39e3095f;
    ram_cell[     386] = 32'h535a8aa9;
    ram_cell[     387] = 32'hc8b5a33b;
    ram_cell[     388] = 32'h0b4067d2;
    ram_cell[     389] = 32'h52004296;
    ram_cell[     390] = 32'h91ec315b;
    ram_cell[     391] = 32'h06ed8685;
    ram_cell[     392] = 32'hffd218e9;
    ram_cell[     393] = 32'h8d286b7a;
    ram_cell[     394] = 32'hfbab2f07;
    ram_cell[     395] = 32'he019e4ac;
    ram_cell[     396] = 32'h2dbd901f;
    ram_cell[     397] = 32'hf6ee9d7e;
    ram_cell[     398] = 32'hb3b02a31;
    ram_cell[     399] = 32'h373c0fce;
    ram_cell[     400] = 32'ha551a874;
    ram_cell[     401] = 32'h4592b1b0;
    ram_cell[     402] = 32'hab3ee921;
    ram_cell[     403] = 32'h4794130c;
    ram_cell[     404] = 32'h5e0e89d8;
    ram_cell[     405] = 32'hc13c1928;
    ram_cell[     406] = 32'h3fc31b64;
    ram_cell[     407] = 32'hec5e531e;
    ram_cell[     408] = 32'hf32cbcb5;
    ram_cell[     409] = 32'h323d9162;
    ram_cell[     410] = 32'h64762c41;
    ram_cell[     411] = 32'h72027e1c;
    ram_cell[     412] = 32'h54cafc94;
    ram_cell[     413] = 32'hc29d0e1c;
    ram_cell[     414] = 32'h460c5caa;
    ram_cell[     415] = 32'h86f5f371;
    ram_cell[     416] = 32'h14feecb5;
    ram_cell[     417] = 32'h23d5e8a1;
    ram_cell[     418] = 32'h33dcf0e4;
    ram_cell[     419] = 32'h1e8bf431;
    ram_cell[     420] = 32'hb294a1cb;
    ram_cell[     421] = 32'h7270f418;
    ram_cell[     422] = 32'hcf51b16f;
    ram_cell[     423] = 32'h3f4531e6;
    ram_cell[     424] = 32'h03d59911;
    ram_cell[     425] = 32'h0007ae86;
    ram_cell[     426] = 32'h45e63a78;
    ram_cell[     427] = 32'haab4e2c7;
    ram_cell[     428] = 32'h319c7db3;
    ram_cell[     429] = 32'h49ee8951;
    ram_cell[     430] = 32'h8c7c9a42;
    ram_cell[     431] = 32'h10d43ab0;
    ram_cell[     432] = 32'he7a04403;
    ram_cell[     433] = 32'h5fab7387;
    ram_cell[     434] = 32'h9ba1f4b6;
    ram_cell[     435] = 32'hdc9cfd5f;
    ram_cell[     436] = 32'h3bd2f963;
    ram_cell[     437] = 32'h84c1c07f;
    ram_cell[     438] = 32'h93e742a7;
    ram_cell[     439] = 32'h476c38ed;
    ram_cell[     440] = 32'h7c590bed;
    ram_cell[     441] = 32'h311e97ed;
    ram_cell[     442] = 32'hc6baa50f;
    ram_cell[     443] = 32'h94eb9033;
    ram_cell[     444] = 32'h51e42933;
    ram_cell[     445] = 32'hb6da1e3d;
    ram_cell[     446] = 32'h40433daf;
    ram_cell[     447] = 32'hfc4d6e88;
    ram_cell[     448] = 32'h4d07eae1;
    ram_cell[     449] = 32'h5ffde31c;
    ram_cell[     450] = 32'hd3f8f6c1;
    ram_cell[     451] = 32'h09e295c9;
    ram_cell[     452] = 32'hd7c12b43;
    ram_cell[     453] = 32'h3e8e3cd7;
    ram_cell[     454] = 32'hf948cb16;
    ram_cell[     455] = 32'h28587129;
    ram_cell[     456] = 32'h64dcad02;
    ram_cell[     457] = 32'h477ecacb;
    ram_cell[     458] = 32'h9c324ac7;
    ram_cell[     459] = 32'h200bf467;
    ram_cell[     460] = 32'h0a8c6792;
    ram_cell[     461] = 32'h4985086e;
    ram_cell[     462] = 32'hca456d80;
    ram_cell[     463] = 32'hb2b2b203;
    ram_cell[     464] = 32'h30506a95;
    ram_cell[     465] = 32'hcb0a035d;
    ram_cell[     466] = 32'hbf23f818;
    ram_cell[     467] = 32'hed9b8e20;
    ram_cell[     468] = 32'h2199dfe6;
    ram_cell[     469] = 32'h8c85b0d6;
    ram_cell[     470] = 32'h1fb73629;
    ram_cell[     471] = 32'h0d8e1021;
    ram_cell[     472] = 32'h2b3e5636;
    ram_cell[     473] = 32'h164c1498;
    ram_cell[     474] = 32'h1f2eadc4;
    ram_cell[     475] = 32'h1c97b73f;
    ram_cell[     476] = 32'h1fb2ef74;
    ram_cell[     477] = 32'h859d6f6b;
    ram_cell[     478] = 32'h7e8d6b0f;
    ram_cell[     479] = 32'hb00b3afc;
    ram_cell[     480] = 32'h66ecdbb0;
    ram_cell[     481] = 32'hc35e8bb3;
    ram_cell[     482] = 32'hd4d0678a;
    ram_cell[     483] = 32'h67f49386;
    ram_cell[     484] = 32'h028912f7;
    ram_cell[     485] = 32'h1ee8f73a;
    ram_cell[     486] = 32'h5f9f06d6;
    ram_cell[     487] = 32'h91993041;
    ram_cell[     488] = 32'h63175aeb;
    ram_cell[     489] = 32'h111409c5;
    ram_cell[     490] = 32'h4d7696fe;
    ram_cell[     491] = 32'ha364c597;
    ram_cell[     492] = 32'hae990aa9;
    ram_cell[     493] = 32'h9d5196af;
    ram_cell[     494] = 32'hb2485967;
    ram_cell[     495] = 32'h0b1730e7;
    ram_cell[     496] = 32'h4c99f17c;
    ram_cell[     497] = 32'hcbe4ff9a;
    ram_cell[     498] = 32'h57b74b0b;
    ram_cell[     499] = 32'hc685c6e2;
    ram_cell[     500] = 32'h502e74f2;
    ram_cell[     501] = 32'hc97fd0da;
    ram_cell[     502] = 32'hd96e2b42;
    ram_cell[     503] = 32'h814732c7;
    ram_cell[     504] = 32'h4e8a36a7;
    ram_cell[     505] = 32'he063c129;
    ram_cell[     506] = 32'h6a5defcf;
    ram_cell[     507] = 32'hd912184f;
    ram_cell[     508] = 32'hcbcc355b;
    ram_cell[     509] = 32'h01b9fad0;
    ram_cell[     510] = 32'h77036ba9;
    ram_cell[     511] = 32'he76e0287;
    // src matrix B
    ram_cell[     512] = 32'hdbde6987;
    ram_cell[     513] = 32'hef86afd7;
    ram_cell[     514] = 32'h39fdb5fc;
    ram_cell[     515] = 32'h3c3a6bb5;
    ram_cell[     516] = 32'he1d4fde9;
    ram_cell[     517] = 32'he57ebe2b;
    ram_cell[     518] = 32'h0f66c56b;
    ram_cell[     519] = 32'h29bef379;
    ram_cell[     520] = 32'h1e8023b7;
    ram_cell[     521] = 32'hf0fda3c9;
    ram_cell[     522] = 32'h8aef1f51;
    ram_cell[     523] = 32'he74bbe55;
    ram_cell[     524] = 32'h6c1822c0;
    ram_cell[     525] = 32'h6505bce2;
    ram_cell[     526] = 32'hfd5ea920;
    ram_cell[     527] = 32'h0a8609ec;
    ram_cell[     528] = 32'h128b00d3;
    ram_cell[     529] = 32'hdbc8ec57;
    ram_cell[     530] = 32'h63f8001b;
    ram_cell[     531] = 32'h0257fbac;
    ram_cell[     532] = 32'hc1e1311b;
    ram_cell[     533] = 32'h6072add0;
    ram_cell[     534] = 32'h0a98ac37;
    ram_cell[     535] = 32'hcb79ecbd;
    ram_cell[     536] = 32'ha749a529;
    ram_cell[     537] = 32'hd255f8a2;
    ram_cell[     538] = 32'h6ad478a5;
    ram_cell[     539] = 32'h3a05d00d;
    ram_cell[     540] = 32'hc1aa0126;
    ram_cell[     541] = 32'h198b587e;
    ram_cell[     542] = 32'heb518f13;
    ram_cell[     543] = 32'h1e074b64;
    ram_cell[     544] = 32'h8986c2fd;
    ram_cell[     545] = 32'h64011af0;
    ram_cell[     546] = 32'h08f80a64;
    ram_cell[     547] = 32'hb646cf50;
    ram_cell[     548] = 32'h2ca257bd;
    ram_cell[     549] = 32'h46d71f72;
    ram_cell[     550] = 32'h684a85ec;
    ram_cell[     551] = 32'hf5a94270;
    ram_cell[     552] = 32'h9eece2be;
    ram_cell[     553] = 32'h486cd751;
    ram_cell[     554] = 32'haaf9eef0;
    ram_cell[     555] = 32'hed43300f;
    ram_cell[     556] = 32'h5db4eafa;
    ram_cell[     557] = 32'hf4d06699;
    ram_cell[     558] = 32'h7e01eb52;
    ram_cell[     559] = 32'h3d3f9614;
    ram_cell[     560] = 32'h8a4a6cd6;
    ram_cell[     561] = 32'hc4d5a0c3;
    ram_cell[     562] = 32'h68b306c1;
    ram_cell[     563] = 32'h65da5755;
    ram_cell[     564] = 32'h206e43d3;
    ram_cell[     565] = 32'h90b51059;
    ram_cell[     566] = 32'h8473ed4f;
    ram_cell[     567] = 32'h1127ac0b;
    ram_cell[     568] = 32'h78c26606;
    ram_cell[     569] = 32'h1617cb04;
    ram_cell[     570] = 32'h7a51087b;
    ram_cell[     571] = 32'h16a0a602;
    ram_cell[     572] = 32'h0d1fbb56;
    ram_cell[     573] = 32'hb05c2e94;
    ram_cell[     574] = 32'h2b840e84;
    ram_cell[     575] = 32'hb70040a4;
    ram_cell[     576] = 32'hb44ddb28;
    ram_cell[     577] = 32'h9ec53126;
    ram_cell[     578] = 32'h1b0fa69f;
    ram_cell[     579] = 32'h836eff23;
    ram_cell[     580] = 32'he4b726e2;
    ram_cell[     581] = 32'h8aefc7ee;
    ram_cell[     582] = 32'haedb7d8e;
    ram_cell[     583] = 32'h245153f6;
    ram_cell[     584] = 32'h6a0694b4;
    ram_cell[     585] = 32'h075f283e;
    ram_cell[     586] = 32'h5f1ee40d;
    ram_cell[     587] = 32'hc4f4fe84;
    ram_cell[     588] = 32'h3dd6f237;
    ram_cell[     589] = 32'h1e7c21f1;
    ram_cell[     590] = 32'h2157e516;
    ram_cell[     591] = 32'h594af9a2;
    ram_cell[     592] = 32'h85ece850;
    ram_cell[     593] = 32'hc36df900;
    ram_cell[     594] = 32'h91254112;
    ram_cell[     595] = 32'h1462ba94;
    ram_cell[     596] = 32'hdf1f57fa;
    ram_cell[     597] = 32'h72050557;
    ram_cell[     598] = 32'had272be0;
    ram_cell[     599] = 32'h7e349054;
    ram_cell[     600] = 32'h2fef861f;
    ram_cell[     601] = 32'h038e54d3;
    ram_cell[     602] = 32'h36d39c30;
    ram_cell[     603] = 32'h039f82e9;
    ram_cell[     604] = 32'hc5bcfbfc;
    ram_cell[     605] = 32'h420f1404;
    ram_cell[     606] = 32'hc4815e60;
    ram_cell[     607] = 32'h9b1f168f;
    ram_cell[     608] = 32'hb8195e5a;
    ram_cell[     609] = 32'hb56f6ee8;
    ram_cell[     610] = 32'ha3062803;
    ram_cell[     611] = 32'hb817d42e;
    ram_cell[     612] = 32'hbc37912e;
    ram_cell[     613] = 32'h8e67005a;
    ram_cell[     614] = 32'h99e62faf;
    ram_cell[     615] = 32'h89f44a70;
    ram_cell[     616] = 32'h6a1a14de;
    ram_cell[     617] = 32'h5638ed8a;
    ram_cell[     618] = 32'h72d68ef5;
    ram_cell[     619] = 32'h72d832ca;
    ram_cell[     620] = 32'hee27ca06;
    ram_cell[     621] = 32'h8d6b4b1c;
    ram_cell[     622] = 32'h883495e5;
    ram_cell[     623] = 32'hde1e372b;
    ram_cell[     624] = 32'h1f3b0b95;
    ram_cell[     625] = 32'h0c5b6895;
    ram_cell[     626] = 32'h275f493c;
    ram_cell[     627] = 32'h6925e41c;
    ram_cell[     628] = 32'hb377c977;
    ram_cell[     629] = 32'hdb1f380a;
    ram_cell[     630] = 32'hf30e304d;
    ram_cell[     631] = 32'h9a786f12;
    ram_cell[     632] = 32'hc85f2b3f;
    ram_cell[     633] = 32'h83338c4b;
    ram_cell[     634] = 32'hd3e56b5e;
    ram_cell[     635] = 32'h27a57cef;
    ram_cell[     636] = 32'h235e0510;
    ram_cell[     637] = 32'ha730aa51;
    ram_cell[     638] = 32'he2fd9d1b;
    ram_cell[     639] = 32'h6d2f3b3e;
    ram_cell[     640] = 32'h1ff60170;
    ram_cell[     641] = 32'h5df88f45;
    ram_cell[     642] = 32'h97ef12cf;
    ram_cell[     643] = 32'h17c4bc75;
    ram_cell[     644] = 32'hb829c33d;
    ram_cell[     645] = 32'h4f65f25b;
    ram_cell[     646] = 32'h674b3ee7;
    ram_cell[     647] = 32'h633d20fb;
    ram_cell[     648] = 32'h661f8f34;
    ram_cell[     649] = 32'h8c33a299;
    ram_cell[     650] = 32'h4a4d4d09;
    ram_cell[     651] = 32'he76f95bc;
    ram_cell[     652] = 32'heae42872;
    ram_cell[     653] = 32'h935f9d89;
    ram_cell[     654] = 32'h7cb653f2;
    ram_cell[     655] = 32'h1d508370;
    ram_cell[     656] = 32'h8ab27955;
    ram_cell[     657] = 32'h6bf27d41;
    ram_cell[     658] = 32'hadc96e3d;
    ram_cell[     659] = 32'h7095808c;
    ram_cell[     660] = 32'h0bf196ff;
    ram_cell[     661] = 32'heeee92c9;
    ram_cell[     662] = 32'haf7fa0da;
    ram_cell[     663] = 32'haaa4c3e2;
    ram_cell[     664] = 32'h68ab81f2;
    ram_cell[     665] = 32'heca69d0c;
    ram_cell[     666] = 32'h29ebca88;
    ram_cell[     667] = 32'h78fff66b;
    ram_cell[     668] = 32'h9c2bc34c;
    ram_cell[     669] = 32'h82b35d83;
    ram_cell[     670] = 32'h39090380;
    ram_cell[     671] = 32'h10bc923e;
    ram_cell[     672] = 32'h4f94bd1d;
    ram_cell[     673] = 32'h974b7507;
    ram_cell[     674] = 32'h61ee5edc;
    ram_cell[     675] = 32'h4573f155;
    ram_cell[     676] = 32'hbec1b512;
    ram_cell[     677] = 32'ha1cb13e4;
    ram_cell[     678] = 32'h7ba2eff9;
    ram_cell[     679] = 32'h2de604e7;
    ram_cell[     680] = 32'he9d68978;
    ram_cell[     681] = 32'h1a5a73d5;
    ram_cell[     682] = 32'h1332c7fb;
    ram_cell[     683] = 32'h98824f65;
    ram_cell[     684] = 32'h2f66bee7;
    ram_cell[     685] = 32'h6cc0ad88;
    ram_cell[     686] = 32'hce21896a;
    ram_cell[     687] = 32'ha436bcd2;
    ram_cell[     688] = 32'h60cd537a;
    ram_cell[     689] = 32'h2341af13;
    ram_cell[     690] = 32'h2657cbc1;
    ram_cell[     691] = 32'h50b821e3;
    ram_cell[     692] = 32'h19f03197;
    ram_cell[     693] = 32'h586c1505;
    ram_cell[     694] = 32'h1b4993ee;
    ram_cell[     695] = 32'h999bc988;
    ram_cell[     696] = 32'h208c231d;
    ram_cell[     697] = 32'h737a8c14;
    ram_cell[     698] = 32'he580e81b;
    ram_cell[     699] = 32'h9c893b81;
    ram_cell[     700] = 32'h1f3de54b;
    ram_cell[     701] = 32'hd889af92;
    ram_cell[     702] = 32'h4d187a9b;
    ram_cell[     703] = 32'h4d816bd2;
    ram_cell[     704] = 32'h55fa7b70;
    ram_cell[     705] = 32'h223fd985;
    ram_cell[     706] = 32'h1e8d3e81;
    ram_cell[     707] = 32'h13a3f9f6;
    ram_cell[     708] = 32'hadfdf58b;
    ram_cell[     709] = 32'h4c97fef7;
    ram_cell[     710] = 32'h703911b6;
    ram_cell[     711] = 32'h76c38552;
    ram_cell[     712] = 32'hd3ab63a7;
    ram_cell[     713] = 32'h7514c536;
    ram_cell[     714] = 32'h26fb77b4;
    ram_cell[     715] = 32'hc3d09010;
    ram_cell[     716] = 32'hd38396b5;
    ram_cell[     717] = 32'h672cedfc;
    ram_cell[     718] = 32'hb9b19743;
    ram_cell[     719] = 32'h20bbf966;
    ram_cell[     720] = 32'hcce4400a;
    ram_cell[     721] = 32'h79ad3471;
    ram_cell[     722] = 32'h73dfa87d;
    ram_cell[     723] = 32'h689de446;
    ram_cell[     724] = 32'h61ae8266;
    ram_cell[     725] = 32'h79247889;
    ram_cell[     726] = 32'h2ed7b8cf;
    ram_cell[     727] = 32'h844e8b5c;
    ram_cell[     728] = 32'h3121fb2d;
    ram_cell[     729] = 32'hc396b79d;
    ram_cell[     730] = 32'h33b74304;
    ram_cell[     731] = 32'h83d89df0;
    ram_cell[     732] = 32'h0e14b6f4;
    ram_cell[     733] = 32'hcec3c5a9;
    ram_cell[     734] = 32'h6f81a454;
    ram_cell[     735] = 32'h8f57cb8a;
    ram_cell[     736] = 32'h7e4e69cc;
    ram_cell[     737] = 32'he33d0441;
    ram_cell[     738] = 32'h6cbeffde;
    ram_cell[     739] = 32'h01113659;
    ram_cell[     740] = 32'h80182562;
    ram_cell[     741] = 32'h7ba669d3;
    ram_cell[     742] = 32'h6c756526;
    ram_cell[     743] = 32'hc6d31742;
    ram_cell[     744] = 32'h60051191;
    ram_cell[     745] = 32'h3da24800;
    ram_cell[     746] = 32'hec16639d;
    ram_cell[     747] = 32'hc09f304c;
    ram_cell[     748] = 32'h4ec4a693;
    ram_cell[     749] = 32'h18950c39;
    ram_cell[     750] = 32'heabb2a46;
    ram_cell[     751] = 32'hb1609c1a;
    ram_cell[     752] = 32'hddb8fd01;
    ram_cell[     753] = 32'h76d7c0fa;
    ram_cell[     754] = 32'h9b64b572;
    ram_cell[     755] = 32'hb6092d4f;
    ram_cell[     756] = 32'h59ce4bc6;
    ram_cell[     757] = 32'h453a7f3f;
    ram_cell[     758] = 32'h35469569;
    ram_cell[     759] = 32'h305cbc95;
    ram_cell[     760] = 32'h53c56f78;
    ram_cell[     761] = 32'h8d40c8f3;
    ram_cell[     762] = 32'h93d8bae4;
    ram_cell[     763] = 32'h0eb9510f;
    ram_cell[     764] = 32'h6fbd49ff;
    ram_cell[     765] = 32'h421f0c7f;
    ram_cell[     766] = 32'h24caedbc;
    ram_cell[     767] = 32'h57509448;
end

endmodule

